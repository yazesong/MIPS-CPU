`timescale 1ns / 1ps

// ��������������ƽ̨
// ֻ���� interface ���裬������ CPU
module tb_peripherals;

  // ʱ�Ӻ͸�λ
  reg clk;
  reg rst;
  
  // �������� IO
  reg  [23:0] switches_in;      // ���뿪������
  wire [7:0]  led_RLD_out;      // ���
  wire [7:0]  led_YLD_out;      // �Ƶ�  
  wire [7:0]  led_GLD_out;      // �̵�
  wire [7:0]  digits_sel_out;   // �����λѡ
  wire [7:0]  digits_data_out;  // ����ܶ�ѡ
  wire        beep_out;         // ������
  reg  [3:0]  keyboard_cols_in; // ����������
  wire [3:0]  keyboard_rows_out;// ���������

  // �����źţ������������裩
  reg  [31:0] bus_addr;
  reg  [31:0] bus_write_data;
  reg         bus_en;
  reg         bus_we;
  reg  [3:0]  bus_byte_sel;
  
  // ������������
  wire [31:0] leds_data_out;
  wire [31:0] switches_data_out;
  wire [31:0] digits_data_out_read;
  wire [31:0] beep_data_out;
  wire [31:0] keyboard_data_out;

  // ʱ������ - 50MHz (20ns period)
  always #10 clk = ~clk;

  // ================================
  // ������������ģ��
  // ================================

  // LED ����
  leds u_leds (
    .rst(rst),
    .clk(clk),
    .addr(bus_addr),
    .en(bus_en),
    .byte_sel(bus_byte_sel),
    .data_in(bus_write_data),
    .we(bus_we),
    .data_out(leds_data_out),
    .RLD(led_RLD_out),
    .YLD(led_YLD_out),
    .GLD(led_GLD_out)
  );

  // ���뿪������
  switches u_switches (
    .rst(rst),
    .clk(clk),
    .addr(bus_addr),
    .en(bus_en),
    .byte_sel(bus_byte_sel),
    .data_in(bus_write_data),
    .we(bus_we),
    .data_out(switches_data_out),
    .switch_in(switches_in)
  );

  // ���������
  digits u_digits (
    .rst(rst),
    .clk(clk),
    .addr(bus_addr),
    .en(bus_en),
    .byte_sel(bus_byte_sel),
    .data_in(bus_write_data),
    .we(bus_we),
    .data_out(digits_data_out_read),
    .sel_out(digits_sel_out),
    .digital_out(digits_data_out)
  );

  // ����������
  beep u_beep (
    .rst(rst),
    .clk(clk),
    .addr(bus_addr),
    .en(bus_en),
    .byte_sel(bus_byte_sel),
    .data_in(bus_write_data),
    .we(bus_we),
    .data_out(beep_data_out),
    .signal_out(beep_out)
  );

  // ��������
  keyboard u_keyboard (
    .rst(rst),
    .clk(clk),
    .addr(bus_addr),
    .en(bus_en),
    .byte_sel(bus_byte_sel),
    .data_in(bus_write_data),
    .we(bus_we),
    .data_out(keyboard_data_out),
    .cols(keyboard_cols_in),
    .rows(keyboard_rows_out)
  );

  // ================================
  // ����������
  // ================================
  initial begin
    // ���� VCD �����ļ�
    $dumpfile("peripherals_waveform.vcd");
    $dumpvars(0, tb_peripherals);
    
    $display("=== ��ʼ�������������� ===");
    
    // ��ʼ��
    clk = 0;
    rst = 1;
    switches_in = 24'h000000;
    keyboard_cols_in = 4'b1111;
    bus_en = 0;
    bus_we = 0;
    bus_addr = 0;
    bus_write_data = 0;
    bus_byte_sel = 4'b1111;
    
    #100;
    rst = 0;
    #100;
    
    // ===================================
    // ���� 1: LED ���� (��ַ: 0xFFFFFC60)
    // ===================================
    $display("���� 1: LED ����");
    bus_addr = 32'hfffffc60;
    bus_write_data = 32'hAABBCCDD;  // R=0xAA, Y=0xBB, G=0xCC
    bus_en = 1;
    bus_we = 1;
    
    #20;  // һ��ʱ������
    
    bus_en = 0;
    bus_we = 0;
    
    $display("LED ��� - R:%h Y:%h G:%h", 
             led_RLD_out, led_YLD_out, led_GLD_out);
    #200;
    
    // ===================================
    // ���� 2: ��ȡ���뿪�� (��ַ: 0xFFFFFC70)
    // ===================================
    $display("���� 2: ���뿪�ض�ȡ");
    switches_in = 24'h123456;  // ���ÿ���ֵ
    
    #100;  // �ȴ�����ֵ������
    
    bus_addr = 32'hfffffc70;
    bus_en = 1;
    bus_we = 0;  // ������
    
    #20;
    
    bus_en = 0;
    
    $display("���ض�ȡֵ: %h", switches_data_out);
    #200;
    
    // ===================================
    // ���� 3: �������ʾ (��ַ: 0xFFFFFC00, 0xFFFFFC04)
    // ===================================
    $display("���� 3: �������ʾ");
    
    // ������ʾ���� (���� 5)
    bus_addr = 32'hfffffc00;
    bus_write_data = 32'd5;
    bus_en = 1;
    bus_we = 1;
    #20;
    bus_en = 0;
    bus_we = 0;
    
    // ����λѡ (�� 0 λ)
    bus_addr = 32'hfffffc04;
    bus_write_data = 32'd0;
    bus_en = 1;
    bus_we = 1;
    #20;
    bus_en = 0;
    bus_we = 0;
    
    $display("����� - λѡ:%h ��ѡ:%h", digits_sel_out, digits_data_out);
    #200;
    
    // ===================================
    // ���� 4: ���������� (��ַ: 0xFFFFFD10)
    // ===================================
    $display("���� 4: ����������");
    
    // �򿪷�����
    bus_addr = 32'hfffffd10;
    bus_write_data = 32'd1;
    bus_en = 1;
    bus_we = 1;
    #20;
    bus_en = 0;
    bus_we = 0;
    
    $display("������״̬ (1=��): %b", beep_out);
    #100;
    
    // �رշ�����
    bus_addr = 32'hfffffd10;
    bus_write_data = 32'd0;
    bus_en = 1;
    bus_we = 1;
    #20;
    bus_en = 0;
    bus_we = 0;
    
    $display("������״̬ (0=��): %b", beep_out);
    #200;
    
    // ===================================
    // ���� 5: ����ɨ�� (�򻯲���)
    // ===================================
    $display("���� 5: ����ɨ�� (��)");
    keyboard_cols_in = 4'b1110;  // ģ�ⰴ������
    
    #500;  // �ȴ�����״̬������
    
    $display("���̶�ȡֵ: %h", keyboard_data_out);
    #200;
    
    // ===================================
    // ��������
    // ===================================
    $display("=== ������������� ===");
    #1000;
    $finish;
  end

endmodule
